module uy(counter1,counter2,counter3,counter4,counter5,counter6,counter7,counter8,control,control2,control3,control4,display,display2,display3,display4,clk,reset,s1,s2,s3,s4,s5,s6,s7,s8,s9);
input clk,reset,s1,s2,s3,s4,s5,s6,s7,s8,s9;
output reg [3:0]control;
output reg [3:0]control2;
output reg [3:0]control3;
output reg [3:0]control4;
output reg [7:0]display;
output reg [7:0]display2;
output reg [7:0]display3;
output reg [7:0]display4;
output reg [3:0]counter1;
output reg [3:0]counter2;
output reg [3:0]counter3;
output reg [3:0]counter4;
output reg [3:0]counter5;
output reg [4:0]counter6;
output reg [4:0]counter7;
output reg [4:0]counter8;
reg clkms,flag1,flag2,clkrms,flag3,flag4;
integer temp1,temp2;
initial
begin
clkms=1'b0;
flag1=1'b0;
flag2=1'b0;
flag3=1'b0;
flag4=1'b0;
temp1=0;
temp2=0;
counter1=4'b0000;
counter2=4'b0000;
counter3=4'b0000;
counter4=4'b0000;
counter5=4'b0000;
counter6=5'b00000;
counter7=5'b00000;
counter8=5'b00000;
end
always@(posedge clk)
begin
temp1=temp1+1;
if(temp1==2000000)
begin
clkms=~clkms;
temp1=0;
end
if(temp2==4000000)
begin
clkrms=~clkrms;
temp2=0;
end
end
always@(posedge clkms)
begin
if(reset==1'b1)
begin
counter1=4'd0;
counter2=4'd0;
counter3=4'd0;
counter4=4'd0;
counter5=5'd0;
counter6=5'd0;
counter7=5'd0;
counter8=5'd0;
end
else if(s1==1'b1)
begin
begin
counter1=counter1+1;
counter2=counter2+1;
counter3=counter3+1;
counter4=counter4+1;
counter5=counter5+1;
counter6=counter6+1;
counter7=counter7+1;
counter8=counter8+1;
end
if(counter1==4'b0001 && s2==1'b1)
begin
flag1=1'b1;
flag2=1'b0;
flag3=1'b0;
flag4=1'b0;
counter2=4'b0000;
counter3=4'b0000;
counter4=4'b0000;
end
else if(counter2==4'b0001 && s3==1'b1)
begin
flag1=1'b0;
flag2=1'b1;
flag3=1'b0;
flag4=1'b0;
counter3=4'b0000;
counter1=4'b0000;
counter4=4'b0000;
end
else if(counter3==4'b0001 && s4==1'b1)
begin
counter1=4'b0000;
counter4=4'b0000;
counter2=4'b0000;
flag1=1'b0;
flag2=1'b0;
flag3=1'b1;
flag4=1'b0;
end
else if(counter4==4'b0001 && s5==1'b1)
begin
counter1=4'b0000;
counter2=4'b0000;
counter3=4'b0000;
flag1=1'b0;
flag2=1'b0;
flag3=1'b0;
flag4=1'b1;
end
else if(counter1 > 4'b0100)
begin
flag1=1'b0;
flag2=1'b0;
flag3=1'b0;
flag4=1'b0;
counter1=4'b0000;
counter2=4'b0000;
counter3=4'b0000;
counter4=4'b0000;
end
else if(s6==1'b1 && counter5 < 4'b1010)
begin
case(counter5)
4'd0: begin
control=4'b0111;
display=8'b11111100;
end
4'd1:begin
control=4'b0111;
display=8'b01100000;
end
4'd2:begin
control=4'b1011;
display=8'b11011010;
end
4'd3:begin
control=4'b1101;
display=8'b11110010;
end
4'd4:begin
control=4'b1110;
display=8'b01100110;
end
4'd5: begin
control=4'b1110;
display=8'b01100110;
end
4'd6:begin
control=4'b1101;
display=8'b11110010;
end
4'd7:begin
control=4'b1011;
display=8'b11011010;
end
4'd8:begin
control=4'b0111;
display=8'b01100000;
end
endcase
end
else if(s7==1'b1 && counter6 < 5'b10010)
begin
case(counter6)
5'd0:begin
control=4'b0111;
display=8'b00000010;
end
5'd1:begin
control=4'b0111;
display=8'b00000010;
end
5'd2:begin
control=4'b1011;
display=8'b00000010;
end
5'd3:begin
control=4'b1101;
display=8'b00000010;
end
5'd4:begin
control=4'b1110;
display=8'b00000010;
end
5'd5:begin
control=4'b1111;
control2=4'b0111;
display2=8'b00000010;
end
5'd6:begin
control=4'b1111;
control2=4'b1011;
display2=8'b00000010;
end
5'd7:begin
control=4'b1111;
control2=4'b1101;
display2=8'b00000010;
end
5'd8:begin
control=4'b1111;
control2=4'b1110;
display2=8'b00000010;
end
5'd9:begin
control=4'b1111;
control2=4'b1111;
control3=4'b0111;
display3=8'b00000010;
end
5'd10:begin
control=4'b1111;
control2=4'b1111;
control3=4'b1011;
display3=8'b00000010;
end
5'd11:begin
control=4'b1111;
control2=4'b1111;
control3=4'b1101;
display3=8'b00000010;
end
5'd12:begin
control=4'b1111;
control2=4'b1111;
control3=4'b1110;
display3=8'b00000010;
end
5'd13:begin
control=4'b1111;
control2=4'b1111;
control3=4'b1111;
control4=4'b0111;
display4=8'b00000010;
end
5'd14:begin
control=4'b1111;
control2=4'b1111;
control3=4'b1111;
control4=4'b1011;
display4=8'b00000010;
end
5'd15:begin
control=4'b1111;
control2=4'b1111;
control3=4'b1111;
control4=4'b1101;
display4=8'b00000010;
end
5'd16:begin
control=4'b1111;
control2=4'b1111;
control3=4'b1111;
control4=4'b1110;
display4=8'b00000010;
end
5'd17:begin
control=4'b1111;
control2=4'b1111;
control3=4'b1111;
control4=4'b1111;
display4=8'b00000010;
counter6=5'd0;
end
endcase

end
else if(s8==1'b1 && counter7 < 5'b10010)
begin
case(counter7)
5'd0:begin
control=4'b0111;
display=8'b11000110;
end
5'd1:begin
control=4'b0111;
display=8'b11000110;
end
5'd2:begin
control=4'b1011;
display=8'b00111010;
end
5'd3:begin
control=4'b1101;
display=8'b11000110;
end
5'd4:begin
control=4'b1110;
display=8'b00111010;
end
5'd5:begin
control=4'b1111;
control2=4'b0111;
display2=8'b11000110;
end
5'd6:begin
control=4'b1111;
control2=4'b1011;
display2=8'b00111010;
end
5'd7:begin
control=4'b1111;
control2=4'b1101;
display2=8'b11000110;
end
5'd8:begin
control=4'b1111;
control2=4'b1110;
display2=8'b00111010;
end
5'd9:begin
control=4'b1111;
control2=4'b1111;
control3=4'b0111;
display3=8'b11000110;
end
5'd10:begin
control=4'b1111;
control2=4'b1111;
control3=4'b1011;
display3=8'b00111010;
end
5'd11:begin
control=4'b1111;
control2=4'b1111;
control3=4'b1101;
display3=8'b11000110;
end
5'd12:begin
control=4'b1111;
control2=4'b1111;
control3=4'b1110;
display3=8'b00111010;
end
5'd13:begin
control=4'b1111;
control2=4'b1111;
control3=4'b1111;
control4=4'b0111;
display4=8'b11000110;
end
5'd14:begin
control=4'b1111;
control2=4'b1111;
control3=4'b1111;
control4=4'b1011;
display4=8'b00111010;
end
5'd15:begin
control=4'b1111;
control2=4'b1111;
control3=4'b1111;
control4=4'b1101;
display4=8'b11000110;
end
5'd16:begin
control=4'b1111;
control2=4'b1111;
control3=4'b1111;
control4=4'b1110;
display4=8'b00111010;
end
5'd17:begin
control=4'b1111;
control2=4'b1111;
control3=4'b1111;
control4=4'b1111;
display4=8'b00000010;
counter6=5'd0;
end
endcase
end
else if(s9==1'b1 && counter8 < 5'b10011)
begin
case(counter7)
5'd0:begin
control=4'b0111;
display=8'b00001000;
end
5'd1:begin
control=4'b0111;
display=8'b00001000;
end
5'd2:begin
control=4'b0111;
display=8'b00000100;
end
5'd3:begin
control=4'b0111;
display=8'b10000000;
end
5'd4:begin
control=4'b0111;
display=8'b01000000;
end
5'd5:begin
control=4'b0111;
display=8'b00100000;
end
5'd6:begin
control=4'b1011;
display=8'b00000100;
end
5'd7:begin
control=4'b1011;
display=8'b10000000;
end
5'd8:begin
control=4'b1011;
display=8'b01000000;
end
5'd9:begin
control=4'b1101;
display=8'b00100000;
end
5'd10:begin
control=4'b1101;
display=8'b00000100;
end
5'd11:begin
control=4'b1101;
display=8'b10000000;
end
5'd12:begin
control=4'b1101;
display=8'b01000000;
end
5'd13:begin
control=4'b1101;
display=8'b00100000;
end
5'd14:begin
control=4'b1110;
display=8'b00100000;
end
5'd15:begin
control=4'b1110;
display=8'b00000100;
end
5'd16:begin
control=4'b1110;
display=8'b10000000;
end
5'd17:begin
control=4'b1110;
display=8'b01000000;
end
5'd18:begin
control=4'b1110;
display=8'b00100000;
counter8=4'd0;
end
endcase

end

if(flag1==1'b1 && s1==1'b1 && flag2==1'b0)
begin
control=4'b0111;
case(counter1)
4'd0:display=8'b11101110;
4'd1:display=8'b11111110;
4'd2:display=8'b10011100;
4'd3:display=8'b10011100;
4'd4:display=8'b11111100;
4'd5:display=8'b10011100;
4'd6:display=8'b10001110;
4'd7:display=8'b01101110;
4'd8:display=8'b01100000;
4'd9:display=8'b11111010;
endcase
end
else if(flag2==1'b1 && s1==1'b1 && flag1==1'b0)
begin
control=4'b1011;
case(counter2)
4'd0:display=8'b11101110;
4'd1:display=8'b11111110;
4'd2:display=8'b10011100;
4'd3:display=8'b10011100;
4'd4:display=8'b11111100;
4'd5:display=8'b10011100;
4'd6:display=8'b10001110;
4'd7:display=8'b01101110;
4'd8:display=8'b01100000;
4'd9:display=8'b11111010;
endcase
end
else if(flag3==1'b1 && s1==1'b1 && flag2==1'b0 )
begin
control=4'b1101;
case(counter3)
4'd0:display=8'b11101110;
4'd1:display=8'b11111110;
4'd2:display=8'b10011100;
4'd3:display=8'b10011100;
4'd4:display=8'b11111100;
4'd5:display=8'b10011100;
4'd6:display=8'b10001110;
4'd7:display=8'b01101110;
4'd8:display=8'b01100000;
4'd9:display=8'b11111010;
endcase

end
else if(flag4==1'b1 && s1==1'b1 && flag3==1'b0 )
begin
control=4'b1110;
case(counter4)
4'd0:display=8'b11101110;
4'd1:display=8'b11111110;
4'd2:display=8'b10011100;
4'd3:display=8'b10011100;
4'd4:display=8'b11111100;
4'd5:display=8'b10011100;
4'd6:display=8'b10001110;
4'd7:display=8'b01101110;
4'd8:display=8'b01100000;
4'd9:display=8'b11111010;
endcase
end

end
end
endmodule
